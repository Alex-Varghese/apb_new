`define num_of_txns 5000
